module fpga_top (
    output wire led
);
    assign led = 1'b0;   // ACTIVE-LOW LED TEST
endmodule
